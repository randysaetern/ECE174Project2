// Forwarding Unit 
// Coded by: Randy Saetern
// Forwards data if necessary

module Forwarding ();




endmodule
