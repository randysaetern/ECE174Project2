module regularALU(input [31:0] I1,I2,output[31:0] out);
	assign out = I1+I2;
endmodule
